library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity mymodule is
	Port (
		input1: in STD_LOGIC_VECTOR (3 downto 0);
		output1: out STD_LOGIC_VECTOR (3 downto 0));
end mymodule;

architecture Behavioral of mymodule is

begin

end Behavioral;
